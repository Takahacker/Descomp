library ieee;
use ieee.std_logic_1164.all;

entity logicaDesvio is
  port (
    entrada_JMP: in std_logic;
    entrada_flag : in std_logic;
    entrada_JEQ : in std_logic;
	 entrada_JSR : in std_logic;
	 entrada_RET : in std_logic;
    saida : out std_logic_vector(1 downto 0)
  );
end entity;

architecture comportamento of logicaDesvio is
  begin
    saida(0) <= entrada_JMP or (entrada_JEQ and entrada_flag) or entrada_JSR;
	 saida(1) <= entrada_RET;
end architecture;